// Data memory

module dmem import config_pkg::*; #(
    // parameter integer RamStart = RamStart;
)(
    input bit [DMemAddrWidth-1:0] address
);

endmodule 
