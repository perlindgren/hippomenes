// Data memory
package dmem_pkg;

  typedef enum {
    BYTE,
    HALFWORD,
    WORD
  } dmem_width_t;

endpackage
