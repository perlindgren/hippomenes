

package a_pkg;

  localparam integer unsigned X = 32;

endpackage
