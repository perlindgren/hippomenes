// Program memory
