// Configuration

