// Instruction decoder