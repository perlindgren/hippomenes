// pc mux
package pc_mux_pkg;
  typedef enum {
    NEXT,
    BRANCH
  } state_t;
endpackage


