// Memory
package mem_pkg;

  typedef enum {
    BYTE = 'b00,
    HALFWORD = 'b10,
    WORD = 'b11
  } mem_width_t;

endpackage
