// Data memory
