// Memory
package mem_pkg;

  typedef enum {
    BYTE,
    HALFWORD,
    WORD
  } mem_width_t;

endpackage
